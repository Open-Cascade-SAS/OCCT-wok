-- SCCS		Date: 04/23/95
--		Information: @(#)MS_InstClass.cdl	1.1
-- File:	MS_InstClass.cdl
-- Created:	Wed Jan 30 12:19:55 1995
-- Author:	Christophe LEYNADIER
--		<cle@ilebon>
---Copyright:	 Matra Datavision 1995


class InstClass 
	---Purpose: 

    from 
    	MS 
    inherits Class from MS
    uses 
     	Type                    from MS,
     	Class                   from MS,
     	GenClass                from MS,
	HAsciiString            from TCollection,
	HSequenceOfHAsciiString from TColStd

is
     
    Create(aName: HAsciiString from TCollection; aPackage: HAsciiString from TCollection) 
    	returns mutable InstClass from MS;

    Validity(me; aName: HAsciiString from TCollection; aPackage: HAsciiString from TCollection);
    	    
    InstType(me : mutable; aType: HAsciiString from TCollection; aPackage: HAsciiString from TCollection);
    InstType(me : mutable;  aType: HAsciiString from TCollection);
    InstTypes(me)
    	returns mutable HSequenceOfHAsciiString from TColStd;
    InstType(me : mutable; aType: Type from MS);
    
    BasicInstType(me : mutable;  aType: HAsciiString from TCollection);
    BasicInstTypes(me)
    	returns mutable HSequenceOfHAsciiString from TColStd;
    ---Purpose: manage the inst types save buffer.
    
    RemoveInstType(me : mutable;  aType: HAsciiString from TCollection);
    ResolveInstType(me : mutable; aType: HAsciiString from TCollection; aTypeConv : HAsciiString from TCollection);
    ---Purpose: the type used to instantiates the generic class
       
    GenType(me: mutable; aType: HAsciiString from TCollection);
    GenTypes(me)
    	returns mutable HSequenceOfHAsciiString from TColStd;
    ---Purpose: the type used to instantiates if the class is nested
    --          they are transformed to inst types when the
    --          method "Instantiates" is called

    GenClass(me: mutable; aName: HAsciiString from TCollection);
    GenClass(me: mutable; aName: HAsciiString from TCollection; aPackage: HAsciiString from TCollection);
    GenClass(me)
    	returns mutable HAsciiString from TCollection;
    ---Purpose: the corresponding generic class.     

    NestedStdClass(me: mutable; aClass : HAsciiString from TCollection);
    NestedInsClass(me: mutable; aClass : HAsciiString from TCollection);
    RemoveNestedStdClass(me: mutable; aClass : HAsciiString from TCollection);
    RemoveNestedInsClass(me: mutable; aClass : HAsciiString from TCollection);
    NestedNeuClass(me: mutable; aClass : HAsciiString from TCollection);
    RemoveNestedNeuClass(me: mutable; aClass : HAsciiString from TCollection);
    ---Purpose: the classes generated by instantiation of a generic
    --          class. 
    --          these classes may contains generics types but
    --          the resolution will occur with a call to the
    --          method "Instantiates"
   
    GetNestedStdClassesName(me)
    	returns mutable HSequenceOfHAsciiString from TColStd;
    GetNestedInsClassesName(me)
    	returns mutable HSequenceOfHAsciiString from TColStd;
    GetNestedNeuClassesName(me)
    	returns mutable HSequenceOfHAsciiString from TColStd;
	    	
    Instantiates(me: mutable);
    ---Purpose: First phase of instantiation
    --          Name and types are created in the metaschema
    --          this is a declaration of all types created by the instantiate command.
   
    InstToStd(me : mutable);
    ---Purpose: Second phase of instantiation.
    --          we create full types
    --          the InstClasses are transformed in StdClasses.
    --          All the generic classes used must be in the MetaSchema    

    IsAlreadyDone(me)
    	returns Boolean from Standard;
    AlreadyDone(me : mutable; flag : Boolean from Standard);
    ---Purpose: test or set the flag when the instantiation has been done

    Initialize(me : mutable);
    ---Purpose: Prepare a instclass for a second instantiates pass
 
      
fields

     myGenClass      : HAsciiString            from TCollection;
     myBasicInsType  : HSequenceOfHAsciiString from TColStd;     -- myInstType save buffer
     myInstType      : HSequenceOfHAsciiString from TColStd;     -- because here we add several inst types during instantiation
     myGenType       : HSequenceOfHAsciiString from TColStd;
     myNestStd       : HSequenceOfHAsciiString from TColStd;
     myNestIns       : HSequenceOfHAsciiString from TColStd;
     myNestNeu       : HSequenceOfHAsciiString from TColStd;
     myComment       : HAsciiString            from TCollection; -- Comment to class declaration 
     myInstFlag      : Boolean from Standard;
     
end InstClass from MS;
