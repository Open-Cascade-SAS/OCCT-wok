-- File:	WOKSH.cdl
-- Created:	Tue Aug  1 23:24:23 1995
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1995

executable WOKSH
is
    
    executable woksh 
    uses
       Tcl_Libs as external
    is
    	woksh;
    end;
    
    executable wokprocess 
    uses
       Tcl_Libs as external
    is
    	wokprocess;
    end;

end;
