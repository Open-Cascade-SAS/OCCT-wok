-- File:	WOKTclTools.cdl
-- Created:	Fri Nov 24 13:59:07 1995
-- Author:	Jean GAUTIER
--		<jga@cobrax>
---Copyright:	 Matra Datavision 1995


package WOKTclTools 

	---Purpose: 

uses

    WOKTools,
    TCollection

is

    imported CommandFunction;
    imported PInterp;
    imported ExitHandler;

    imported WokCommand;
    
    class Package;

    class Interpretor;

    generic class HandleTable;

    class MsgAPI;

--    class SequenceOfHandleTable 
--    	instantiates Sequence from TCollection ( HandleTable from WOKTclTools);

end WOKTclTools;
