-- File:	MS_Imported.cdl
-- Created:	Mon Aug 23 18:44:03 1993
-- Author:	Christophe LEYNADIER
--		<cle@ilebon>
---Copyright:	 Matra Datavision 1993

class Imported 
	---Purpose: 

    from 
    	MS 
    inherits NatType from MS
    uses 
    	HSequenceOfHAsciiString from TColStd,
	HAsciiString from TCollection

is

    Create(aName, aPackage, aContainer: HAsciiString; aPrivate: Boolean) 
    	returns mutable Imported from MS;

    IsTransient(me)
    	returns Boolean from Standard;

    SetTransient(me : mutable; theValue : Boolean from Standard) is static;

fields

  myIsTransient : Boolean from Standard;

end Imported from MS;
