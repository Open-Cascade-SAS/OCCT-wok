-- SCCS		Date: 04/23/95
--		Information: @(#)MS_Enum.cdl	1.1
-- File:	MS_Enum.cdl
-- Created:	Wed Jan 30 12:38:17 1995
-- Author:	Christophe LEYNADIER
--		<cle@ilebon>
---Copyright:	 Matra Datavision 1995


class Enum 
	---Purpose: 

    from 
    	MS 
    inherits NatType from MS
    uses 
    	HSequenceOfHAsciiString from TColStd,
	HAsciiString from TCollection

is

    Create(aName, aPackage, aContainer: HAsciiString; aPrivate: Boolean) 
    	returns mutable Enum from MS;
    
    Enum(me: mutable; aEnum: HAsciiString);
    Enums(me)
    	returns mutable HSequenceOfHAsciiString from TColStd;
	
    Check(me);

fields

    myEnums        : HSequenceOfHAsciiString from TColStd;

end Enum from MS;








